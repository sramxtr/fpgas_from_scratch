
module debouncer(
    input logic clk,
    input logic button_in,
    output logic button_out
    );
    
    // TODO
    
endmodule
