
module button_to_led_top(
    input button_in,
    output led_out
    );
    
    assign led_out = button_in;
    
endmodule
