
module rising_edge_to_pulse(
    input logic clk,
    input logic data_in,
    output logic data_out
    );
    
    // TODO
    
endmodule
