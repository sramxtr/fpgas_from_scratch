
module pattern_checker(
    input logic clk,
    input logic reset,
    input logic action_in,
    input logic [3:0] code_in,
    output logic led_r_out,
    output logic led_g_out,
    output logic led_b_out
    );
    
    // TODO
    
endmodule
